module gac_not_gate_6_BHV (x, z);
  input [5:0] x;
  output [5:0] z;
  
  assign z = ~x ;
  
endmodule
  



