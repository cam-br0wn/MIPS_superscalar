module gac_not_gate (x, z);
  input x;
  output z;
  
  assign z = ~x ;
  
  
endmodule
  




