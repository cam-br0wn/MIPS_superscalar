module gac_not_gate_32 (x, z);
  input [31:0] x;
  output [31:0] z;
  
  assign z = ~x ;
  
  
endmodule
  


